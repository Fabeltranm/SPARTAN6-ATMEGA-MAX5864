module sum4bcc (xi, yi, ci,co,zi);

// completar  para que la descripción funciones

  input [3 :0] xi;
  input [3 :0] yi;
  input  ci;
  output co;
  output [3 :0] zi;

  wire c1
  sum1bcc s0(.xi(x[0]), .yi(y[0]), .ci(ci), .co(c1) ,.zi(z[0]));
  // sum1bcc s1 ...
  // sum1bcc s2 ...
  // sum1bcc s3 ...


endmodule
